------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnologa Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=14); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

library synplify;
architecture rtl of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);
   attribute syn_ramstyle : string;
   attribute syn_ramstyle of addr_r : signal is "block_ram";

   signal ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80cfd00c",
     3 => x"3a0b0b80",
     4 => x"c7d80400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80c8a02d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80cf",
   162 => x"bc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8d",
   171 => x"d32d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8f",
   179 => x"852d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80cfcc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81943f80",
   257 => x"c6e23f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"ff3d0d80",
   281 => x"dfbc3351",
   282 => x"70a73880",
   283 => x"cfd80870",
   284 => x"08525270",
   285 => x"802e9438",
   286 => x"841280cf",
   287 => x"d80c702d",
   288 => x"80cfd808",
   289 => x"70085252",
   290 => x"70ee3881",
   291 => x"0b80dfbc",
   292 => x"34833d0d",
   293 => x"0404803d",
   294 => x"0d0b0b80",
   295 => x"dfb40880",
   296 => x"2e8e380b",
   297 => x"0b0b0b80",
   298 => x"0b802e09",
   299 => x"81068538",
   300 => x"823d0d04",
   301 => x"0b0b80df",
   302 => x"b4510b0b",
   303 => x"0bf6c13f",
   304 => x"823d0d04",
   305 => x"04ff3d0d",
   306 => x"0b0b80cf",
   307 => x"945189d8",
   308 => x"3f71800c",
   309 => x"833d0d04",
   310 => x"fe3d0d80",
   311 => x"dfc00853",
   312 => x"84130870",
   313 => x"882a7081",
   314 => x"06515252",
   315 => x"70802ef0",
   316 => x"387181ff",
   317 => x"06800c84",
   318 => x"3d0d04ff",
   319 => x"3d0d80df",
   320 => x"c0085271",
   321 => x"0870882a",
   322 => x"81327081",
   323 => x"06515151",
   324 => x"70f13873",
   325 => x"720c833d",
   326 => x"0d0480cf",
   327 => x"cc08802e",
   328 => x"80c43880",
   329 => x"cfd00882",
   330 => x"2e098106",
   331 => x"9f3880c0",
   332 => x"a9808c0b",
   333 => x"80dfc00c",
   334 => x"80c0a980",
   335 => x"940b80df",
   336 => x"c40c80cf",
   337 => x"a40b80df",
   338 => x"b80cb939",
   339 => x"8380800b",
   340 => x"80dfc00c",
   341 => x"82a0800b",
   342 => x"80dfc40c",
   343 => x"8290800b",
   344 => x"80dfb80c",
   345 => x"9f39f880",
   346 => x"8080a40b",
   347 => x"80dfc00c",
   348 => x"f8808082",
   349 => x"800b80df",
   350 => x"c40cf880",
   351 => x"8084800b",
   352 => x"80dfb80c",
   353 => x"04f33d0d",
   354 => x"7f80dfc4",
   355 => x"08565c82",
   356 => x"750c8059",
   357 => x"805a805b",
   358 => x"7a842980",
   359 => x"dfc40805",
   360 => x"70087108",
   361 => x"719f2c7e",
   362 => x"852b5855",
   363 => x"55913df8",
   364 => x"05535957",
   365 => x"a83f7c7e",
   366 => x"7a72077c",
   367 => x"72077171",
   368 => x"60810541",
   369 => x"5f5d5b59",
   370 => x"5755817b",
   371 => x"27ca3876",
   372 => x"7c0c7784",
   373 => x"1d0c7b80",
   374 => x"0c8f3d0d",
   375 => x"048c0802",
   376 => x"8c0cf53d",
   377 => x"0d8c0894",
   378 => x"05089d38",
   379 => x"8c088c05",
   380 => x"088c0890",
   381 => x"05088c08",
   382 => x"88050858",
   383 => x"56547376",
   384 => x"0c748417",
   385 => x"0c81bf39",
   386 => x"800b8c08",
   387 => x"f0050c80",
   388 => x"0b8c08f4",
   389 => x"050c8c08",
   390 => x"8c05088c",
   391 => x"08900508",
   392 => x"5654738c",
   393 => x"08f0050c",
   394 => x"748c08f4",
   395 => x"050c8c08",
   396 => x"f8058c08",
   397 => x"f0055656",
   398 => x"88705475",
   399 => x"53765254",
   400 => x"858d3fa0",
   401 => x"0b8c0894",
   402 => x"0508318c",
   403 => x"08ec050c",
   404 => x"8c08ec05",
   405 => x"0880249d",
   406 => x"38800b8c",
   407 => x"08f4050c",
   408 => x"8c08ec05",
   409 => x"08308c08",
   410 => x"fc050871",
   411 => x"2b8c08f0",
   412 => x"050c54b9",
   413 => x"398c08fc",
   414 => x"05088c08",
   415 => x"ec05082a",
   416 => x"8c08e805",
   417 => x"0c8c08fc",
   418 => x"05088c08",
   419 => x"9405082b",
   420 => x"8c08f405",
   421 => x"0c8c08f8",
   422 => x"05088c08",
   423 => x"9405082b",
   424 => x"708c08e8",
   425 => x"0508078c",
   426 => x"08f0050c",
   427 => x"548c08f0",
   428 => x"05088c08",
   429 => x"f405088c",
   430 => x"08880508",
   431 => x"58565473",
   432 => x"760c7484",
   433 => x"170c8c08",
   434 => x"88050880",
   435 => x"0c8d3d0d",
   436 => x"8c0c048c",
   437 => x"08028c0c",
   438 => x"f93d0d80",
   439 => x"0b8c08fc",
   440 => x"050c8c08",
   441 => x"88050880",
   442 => x"25ab388c",
   443 => x"08880508",
   444 => x"308c0888",
   445 => x"050c800b",
   446 => x"8c08f405",
   447 => x"0c8c08fc",
   448 => x"05088838",
   449 => x"810b8c08",
   450 => x"f4050c8c",
   451 => x"08f40508",
   452 => x"8c08fc05",
   453 => x"0c8c088c",
   454 => x"05088025",
   455 => x"ab388c08",
   456 => x"8c050830",
   457 => x"8c088c05",
   458 => x"0c800b8c",
   459 => x"08f0050c",
   460 => x"8c08fc05",
   461 => x"08883881",
   462 => x"0b8c08f0",
   463 => x"050c8c08",
   464 => x"f005088c",
   465 => x"08fc050c",
   466 => x"80538c08",
   467 => x"8c050852",
   468 => x"8c088805",
   469 => x"085181a7",
   470 => x"3f800870",
   471 => x"8c08f805",
   472 => x"0c548c08",
   473 => x"fc050880",
   474 => x"2e8c388c",
   475 => x"08f80508",
   476 => x"308c08f8",
   477 => x"050c8c08",
   478 => x"f8050870",
   479 => x"800c5489",
   480 => x"3d0d8c0c",
   481 => x"048c0802",
   482 => x"8c0cfb3d",
   483 => x"0d800b8c",
   484 => x"08fc050c",
   485 => x"8c088805",
   486 => x"08802593",
   487 => x"388c0888",
   488 => x"0508308c",
   489 => x"0888050c",
   490 => x"810b8c08",
   491 => x"fc050c8c",
   492 => x"088c0508",
   493 => x"80258c38",
   494 => x"8c088c05",
   495 => x"08308c08",
   496 => x"8c050c81",
   497 => x"538c088c",
   498 => x"0508528c",
   499 => x"08880508",
   500 => x"51ad3f80",
   501 => x"08708c08",
   502 => x"f8050c54",
   503 => x"8c08fc05",
   504 => x"08802e8c",
   505 => x"388c08f8",
   506 => x"0508308c",
   507 => x"08f8050c",
   508 => x"8c08f805",
   509 => x"0870800c",
   510 => x"54873d0d",
   511 => x"8c0c048c",
   512 => x"08028c0c",
   513 => x"fd3d0d81",
   514 => x"0b8c08fc",
   515 => x"050c800b",
   516 => x"8c08f805",
   517 => x"0c8c088c",
   518 => x"05088c08",
   519 => x"88050827",
   520 => x"ac388c08",
   521 => x"fc050880",
   522 => x"2ea33880",
   523 => x"0b8c088c",
   524 => x"05082499",
   525 => x"388c088c",
   526 => x"0508108c",
   527 => x"088c050c",
   528 => x"8c08fc05",
   529 => x"08108c08",
   530 => x"fc050cc9",
   531 => x"398c08fc",
   532 => x"0508802e",
   533 => x"80c9388c",
   534 => x"088c0508",
   535 => x"8c088805",
   536 => x"0826a138",
   537 => x"8c088805",
   538 => x"088c088c",
   539 => x"0508318c",
   540 => x"0888050c",
   541 => x"8c08f805",
   542 => x"088c08fc",
   543 => x"0508078c",
   544 => x"08f8050c",
   545 => x"8c08fc05",
   546 => x"08812a8c",
   547 => x"08fc050c",
   548 => x"8c088c05",
   549 => x"08812a8c",
   550 => x"088c050c",
   551 => x"ffaf398c",
   552 => x"08900508",
   553 => x"802e8f38",
   554 => x"8c088805",
   555 => x"08708c08",
   556 => x"f4050c51",
   557 => x"8d398c08",
   558 => x"f8050870",
   559 => x"8c08f405",
   560 => x"0c518c08",
   561 => x"f4050880",
   562 => x"0c853d0d",
   563 => x"8c0c04fc",
   564 => x"3d0d7670",
   565 => x"797b5555",
   566 => x"55558f72",
   567 => x"278c3872",
   568 => x"75078306",
   569 => x"5170802e",
   570 => x"a738ff12",
   571 => x"5271ff2e",
   572 => x"98387270",
   573 => x"81055433",
   574 => x"74708105",
   575 => x"5634ff12",
   576 => x"5271ff2e",
   577 => x"098106ea",
   578 => x"3874800c",
   579 => x"863d0d04",
   580 => x"74517270",
   581 => x"84055408",
   582 => x"71708405",
   583 => x"530c7270",
   584 => x"84055408",
   585 => x"71708405",
   586 => x"530c7270",
   587 => x"84055408",
   588 => x"71708405",
   589 => x"530c7270",
   590 => x"84055408",
   591 => x"71708405",
   592 => x"530cf012",
   593 => x"52718f26",
   594 => x"c9388372",
   595 => x"27953872",
   596 => x"70840554",
   597 => x"08717084",
   598 => x"05530cfc",
   599 => x"12527183",
   600 => x"26ed3870",
   601 => x"54ff8339",
   602 => x"f73d0d7c",
   603 => x"70525380",
   604 => x"c83f7254",
   605 => x"80085580",
   606 => x"cfa85681",
   607 => x"57800881",
   608 => x"055a8b3d",
   609 => x"e4115953",
   610 => x"8259f413",
   611 => x"527b8811",
   612 => x"08525381",
   613 => x"833f8008",
   614 => x"30708008",
   615 => x"079f2c8a",
   616 => x"07800c53",
   617 => x"8b3d0d04",
   618 => x"ff3d0d73",
   619 => x"5280cfdc",
   620 => x"0851ffb4",
   621 => x"3f833d0d",
   622 => x"04fd3d0d",
   623 => x"75707183",
   624 => x"06535552",
   625 => x"70b83871",
   626 => x"70087009",
   627 => x"f7fbfdff",
   628 => x"120670f8",
   629 => x"84828180",
   630 => x"06515152",
   631 => x"53709d38",
   632 => x"84137008",
   633 => x"7009f7fb",
   634 => x"fdff1206",
   635 => x"70f88482",
   636 => x"81800651",
   637 => x"51525370",
   638 => x"802ee538",
   639 => x"72527133",
   640 => x"5170802e",
   641 => x"8a388112",
   642 => x"70335252",
   643 => x"70f83871",
   644 => x"7431800c",
   645 => x"853d0d04",
   646 => x"f23d0d60",
   647 => x"62881108",
   648 => x"7057575f",
   649 => x"5a74802e",
   650 => x"8190388c",
   651 => x"1a227083",
   652 => x"2a813270",
   653 => x"81065155",
   654 => x"58738638",
   655 => x"901a0891",
   656 => x"38795190",
   657 => x"a23fff54",
   658 => x"800880ee",
   659 => x"388c1a22",
   660 => x"587d0857",
   661 => x"807883ff",
   662 => x"ff06700a",
   663 => x"100a7081",
   664 => x"06515657",
   665 => x"5573752e",
   666 => x"80d73874",
   667 => x"90387608",
   668 => x"84180888",
   669 => x"19595659",
   670 => x"74802ef2",
   671 => x"38745488",
   672 => x"80752784",
   673 => x"38888054",
   674 => x"73537852",
   675 => x"9c1a0851",
   676 => x"a41a0854",
   677 => x"732d800b",
   678 => x"80082582",
   679 => x"e6388008",
   680 => x"19758008",
   681 => x"317f8805",
   682 => x"08800831",
   683 => x"70618805",
   684 => x"0c565659",
   685 => x"73ffb438",
   686 => x"80547380",
   687 => x"0c903d0d",
   688 => x"04758132",
   689 => x"70810676",
   690 => x"41515473",
   691 => x"802e81c1",
   692 => x"38749038",
   693 => x"76088418",
   694 => x"08881959",
   695 => x"56597480",
   696 => x"2ef23888",
   697 => x"1a087883",
   698 => x"ffff0670",
   699 => x"892a7081",
   700 => x"06515659",
   701 => x"5673802e",
   702 => x"82fa3875",
   703 => x"75278d38",
   704 => x"77872a70",
   705 => x"81065154",
   706 => x"7382b538",
   707 => x"74762783",
   708 => x"38745675",
   709 => x"53785279",
   710 => x"08518582",
   711 => x"3f881a08",
   712 => x"7631881b",
   713 => x"0c790816",
   714 => x"7a0c7456",
   715 => x"75197577",
   716 => x"317f8805",
   717 => x"08783170",
   718 => x"6188050c",
   719 => x"56565973",
   720 => x"802efef4",
   721 => x"388c1a22",
   722 => x"58ff8639",
   723 => x"77785479",
   724 => x"537b5256",
   725 => x"84c83f88",
   726 => x"1a087831",
   727 => x"881b0c79",
   728 => x"08187a0c",
   729 => x"7c76315d",
   730 => x"7c8e3879",
   731 => x"518fdc3f",
   732 => x"8008818f",
   733 => x"3880085f",
   734 => x"75197577",
   735 => x"317f8805",
   736 => x"08783170",
   737 => x"6188050c",
   738 => x"56565973",
   739 => x"802efea8",
   740 => x"38748183",
   741 => x"38760884",
   742 => x"18088819",
   743 => x"59565974",
   744 => x"802ef238",
   745 => x"74538a52",
   746 => x"785182d3",
   747 => x"3f800879",
   748 => x"3181055d",
   749 => x"80088438",
   750 => x"81155d81",
   751 => x"5f7c5874",
   752 => x"7d278338",
   753 => x"7458941a",
   754 => x"08881b08",
   755 => x"11575c80",
   756 => x"7a085c54",
   757 => x"901a087b",
   758 => x"27833881",
   759 => x"54757825",
   760 => x"843873ba",
   761 => x"387b7824",
   762 => x"fee2387b",
   763 => x"5378529c",
   764 => x"1a0851a4",
   765 => x"1a085473",
   766 => x"2d800856",
   767 => x"80088024",
   768 => x"fee2388c",
   769 => x"1a2280c0",
   770 => x"0754738c",
   771 => x"1b23ff54",
   772 => x"73800c90",
   773 => x"3d0d047e",
   774 => x"ffa338ff",
   775 => x"87397553",
   776 => x"78527a51",
   777 => x"82f83f79",
   778 => x"08167a0c",
   779 => x"79518e9b",
   780 => x"3f8008cf",
   781 => x"387c7631",
   782 => x"5d7cfebc",
   783 => x"38feac39",
   784 => x"901a087a",
   785 => x"08713176",
   786 => x"1170565a",
   787 => x"575280cf",
   788 => x"dc085184",
   789 => x"8c3f8008",
   790 => x"802effa7",
   791 => x"38800890",
   792 => x"1b0c8008",
   793 => x"167a0c77",
   794 => x"941b0c74",
   795 => x"881b0c74",
   796 => x"56fd9939",
   797 => x"79085890",
   798 => x"1a087827",
   799 => x"83388154",
   800 => x"75752784",
   801 => x"3873b338",
   802 => x"941a0856",
   803 => x"75752680",
   804 => x"d3387553",
   805 => x"78529c1a",
   806 => x"0851a41a",
   807 => x"0854732d",
   808 => x"80085680",
   809 => x"088024fd",
   810 => x"83388c1a",
   811 => x"2280c007",
   812 => x"54738c1b",
   813 => x"23ff54fe",
   814 => x"d7397553",
   815 => x"78527751",
   816 => x"81dc3f79",
   817 => x"08167a0c",
   818 => x"79518cff",
   819 => x"3f800880",
   820 => x"2efcd938",
   821 => x"8c1a2280",
   822 => x"c0075473",
   823 => x"8c1b23ff",
   824 => x"54fead39",
   825 => x"74755479",
   826 => x"53785256",
   827 => x"81b03f88",
   828 => x"1a087531",
   829 => x"881b0c79",
   830 => x"08157a0c",
   831 => x"fcae39fa",
   832 => x"3d0d7a79",
   833 => x"028805a7",
   834 => x"05335652",
   835 => x"53837327",
   836 => x"8a387083",
   837 => x"06527180",
   838 => x"2ea838ff",
   839 => x"135372ff",
   840 => x"2e973870",
   841 => x"33527372",
   842 => x"2e913881",
   843 => x"11ff1454",
   844 => x"5172ff2e",
   845 => x"098106eb",
   846 => x"38805170",
   847 => x"800c883d",
   848 => x"0d047072",
   849 => x"57558351",
   850 => x"75828029",
   851 => x"14ff1252",
   852 => x"56708025",
   853 => x"f3388373",
   854 => x"27bf3874",
   855 => x"08763270",
   856 => x"09f7fbfd",
   857 => x"ff120670",
   858 => x"f8848281",
   859 => x"80065151",
   860 => x"5170802e",
   861 => x"99387451",
   862 => x"80527033",
   863 => x"5773772e",
   864 => x"ffb93881",
   865 => x"11811353",
   866 => x"51837227",
   867 => x"ed38fc13",
   868 => x"84165653",
   869 => x"728326c3",
   870 => x"387451fe",
   871 => x"fe39fa3d",
   872 => x"0d787a7c",
   873 => x"72727257",
   874 => x"57575956",
   875 => x"56747627",
   876 => x"b2387615",
   877 => x"51757127",
   878 => x"aa387077",
   879 => x"17ff1454",
   880 => x"555371ff",
   881 => x"2e9638ff",
   882 => x"14ff1454",
   883 => x"54723374",
   884 => x"34ff1252",
   885 => x"71ff2e09",
   886 => x"8106ec38",
   887 => x"75800c88",
   888 => x"3d0d0476",
   889 => x"8f269738",
   890 => x"ff125271",
   891 => x"ff2eed38",
   892 => x"72708105",
   893 => x"54337470",
   894 => x"81055634",
   895 => x"eb397476",
   896 => x"07830651",
   897 => x"70e23875",
   898 => x"75545172",
   899 => x"70840554",
   900 => x"08717084",
   901 => x"05530c72",
   902 => x"70840554",
   903 => x"08717084",
   904 => x"05530c72",
   905 => x"70840554",
   906 => x"08717084",
   907 => x"05530c72",
   908 => x"70840554",
   909 => x"08717084",
   910 => x"05530cf0",
   911 => x"1252718f",
   912 => x"26c93883",
   913 => x"72279538",
   914 => x"72708405",
   915 => x"54087170",
   916 => x"8405530c",
   917 => x"fc125271",
   918 => x"8326ed38",
   919 => x"7054ff88",
   920 => x"39ef3d0d",
   921 => x"63656740",
   922 => x"5d427b80",
   923 => x"2e84fa38",
   924 => x"6151a5b6",
   925 => x"3ff81c70",
   926 => x"84120870",
   927 => x"fc067062",
   928 => x"8b0570f8",
   929 => x"06415945",
   930 => x"5b5c4157",
   931 => x"96742782",
   932 => x"c338807b",
   933 => x"247e7c26",
   934 => x"07598054",
   935 => x"78742e09",
   936 => x"810682a9",
   937 => x"38777b25",
   938 => x"81fc3877",
   939 => x"1780d798",
   940 => x"0b880508",
   941 => x"5e567c76",
   942 => x"2e84bd38",
   943 => x"84160870",
   944 => x"fe061784",
   945 => x"11088106",
   946 => x"51555573",
   947 => x"828b3874",
   948 => x"fc06597c",
   949 => x"762e84dd",
   950 => x"3877195f",
   951 => x"7e7b2581",
   952 => x"fd387981",
   953 => x"06547382",
   954 => x"bf387677",
   955 => x"08318411",
   956 => x"08fc0656",
   957 => x"5a75802e",
   958 => x"91387c76",
   959 => x"2e84ea38",
   960 => x"74191859",
   961 => x"787b2584",
   962 => x"89387980",
   963 => x"2e829938",
   964 => x"7715567a",
   965 => x"76248290",
   966 => x"388c1a08",
   967 => x"881b0871",
   968 => x"8c120c88",
   969 => x"120c5579",
   970 => x"76595788",
   971 => x"1761fc05",
   972 => x"575975a4",
   973 => x"2685ef38",
   974 => x"7b795555",
   975 => x"93762780",
   976 => x"c9387b70",
   977 => x"84055d08",
   978 => x"7c56790c",
   979 => x"74708405",
   980 => x"56088c18",
   981 => x"0c901754",
   982 => x"9b7627ae",
   983 => x"38747084",
   984 => x"05560874",
   985 => x"0c747084",
   986 => x"05560894",
   987 => x"180c9817",
   988 => x"54a37627",
   989 => x"95387470",
   990 => x"84055608",
   991 => x"740c7470",
   992 => x"84055608",
   993 => x"9c180ca0",
   994 => x"17547470",
   995 => x"84055608",
   996 => x"74708405",
   997 => x"560c7470",
   998 => x"84055608",
   999 => x"74708405",
  1000 => x"560c7408",
  1001 => x"740c777b",
  1002 => x"3156758f",
  1003 => x"2680c938",
  1004 => x"84170881",
  1005 => x"06780784",
  1006 => x"180c7717",
  1007 => x"84110881",
  1008 => x"0784120c",
  1009 => x"546151a2",
  1010 => x"e23f8817",
  1011 => x"5473800c",
  1012 => x"933d0d04",
  1013 => x"905bfdba",
  1014 => x"397856fe",
  1015 => x"85398c16",
  1016 => x"08881708",
  1017 => x"718c120c",
  1018 => x"88120c55",
  1019 => x"7e707c31",
  1020 => x"57588f76",
  1021 => x"27ffb938",
  1022 => x"7a178418",
  1023 => x"0881067c",
  1024 => x"0784190c",
  1025 => x"76810784",
  1026 => x"120c7611",
  1027 => x"84110881",
  1028 => x"0784120c",
  1029 => x"55880552",
  1030 => x"61518cf7",
  1031 => x"3f6151a2",
  1032 => x"8a3f8817",
  1033 => x"54ffa639",
  1034 => x"7d526151",
  1035 => x"94f73f80",
  1036 => x"08598008",
  1037 => x"802e81a3",
  1038 => x"388008f8",
  1039 => x"05608405",
  1040 => x"08fe0661",
  1041 => x"05555776",
  1042 => x"742e83e6",
  1043 => x"38fc1856",
  1044 => x"75a42681",
  1045 => x"aa387b80",
  1046 => x"08555593",
  1047 => x"762780d8",
  1048 => x"38747084",
  1049 => x"05560880",
  1050 => x"08708405",
  1051 => x"800c0c80",
  1052 => x"08757084",
  1053 => x"05570871",
  1054 => x"70840553",
  1055 => x"0c549b76",
  1056 => x"27b63874",
  1057 => x"70840556",
  1058 => x"08747084",
  1059 => x"05560c74",
  1060 => x"70840556",
  1061 => x"08747084",
  1062 => x"05560ca3",
  1063 => x"76279938",
  1064 => x"74708405",
  1065 => x"56087470",
  1066 => x"8405560c",
  1067 => x"74708405",
  1068 => x"56087470",
  1069 => x"8405560c",
  1070 => x"74708405",
  1071 => x"56087470",
  1072 => x"8405560c",
  1073 => x"74708405",
  1074 => x"56087470",
  1075 => x"8405560c",
  1076 => x"7408740c",
  1077 => x"7b526151",
  1078 => x"8bb93f61",
  1079 => x"51a0cc3f",
  1080 => x"78547380",
  1081 => x"0c933d0d",
  1082 => x"047d5261",
  1083 => x"5193b63f",
  1084 => x"8008800c",
  1085 => x"933d0d04",
  1086 => x"84160855",
  1087 => x"fbd13975",
  1088 => x"537b5280",
  1089 => x"0851efc7",
  1090 => x"3f7b5261",
  1091 => x"518b843f",
  1092 => x"ca398c16",
  1093 => x"08881708",
  1094 => x"718c120c",
  1095 => x"88120c55",
  1096 => x"8c1a0888",
  1097 => x"1b08718c",
  1098 => x"120c8812",
  1099 => x"0c557979",
  1100 => x"5957fbf7",
  1101 => x"39771990",
  1102 => x"1c555573",
  1103 => x"7524fba2",
  1104 => x"387a1770",
  1105 => x"80d7980b",
  1106 => x"88050c75",
  1107 => x"7c318107",
  1108 => x"84120c5d",
  1109 => x"84170881",
  1110 => x"067b0784",
  1111 => x"180c6151",
  1112 => x"9fc93f88",
  1113 => x"1754fce5",
  1114 => x"39741918",
  1115 => x"901c555d",
  1116 => x"737d24fb",
  1117 => x"95388c1a",
  1118 => x"08881b08",
  1119 => x"718c120c",
  1120 => x"88120c55",
  1121 => x"881a61fc",
  1122 => x"05575975",
  1123 => x"a42681ae",
  1124 => x"387b7955",
  1125 => x"55937627",
  1126 => x"80c9387b",
  1127 => x"7084055d",
  1128 => x"087c5679",
  1129 => x"0c747084",
  1130 => x"0556088c",
  1131 => x"1b0c901a",
  1132 => x"549b7627",
  1133 => x"ae387470",
  1134 => x"84055608",
  1135 => x"740c7470",
  1136 => x"84055608",
  1137 => x"941b0c98",
  1138 => x"1a54a376",
  1139 => x"27953874",
  1140 => x"70840556",
  1141 => x"08740c74",
  1142 => x"70840556",
  1143 => x"089c1b0c",
  1144 => x"a01a5474",
  1145 => x"70840556",
  1146 => x"08747084",
  1147 => x"05560c74",
  1148 => x"70840556",
  1149 => x"08747084",
  1150 => x"05560c74",
  1151 => x"08740c7a",
  1152 => x"1a7080d7",
  1153 => x"980b8805",
  1154 => x"0c7d7c31",
  1155 => x"81078412",
  1156 => x"0c54841a",
  1157 => x"0881067b",
  1158 => x"07841b0c",
  1159 => x"61519e8b",
  1160 => x"3f7854fd",
  1161 => x"bd397553",
  1162 => x"7b527851",
  1163 => x"eda13ffa",
  1164 => x"f5398417",
  1165 => x"08fc0618",
  1166 => x"605858fa",
  1167 => x"e9397553",
  1168 => x"7b527851",
  1169 => x"ed893f7a",
  1170 => x"1a7080d7",
  1171 => x"980b8805",
  1172 => x"0c7d7c31",
  1173 => x"81078412",
  1174 => x"0c54841a",
  1175 => x"0881067b",
  1176 => x"07841b0c",
  1177 => x"ffb639fa",
  1178 => x"3d0d7880",
  1179 => x"cfdc0854",
  1180 => x"55b81308",
  1181 => x"802e81b6",
  1182 => x"388c1522",
  1183 => x"7083ffff",
  1184 => x"0670832a",
  1185 => x"81327081",
  1186 => x"06515555",
  1187 => x"5672802e",
  1188 => x"80dc3873",
  1189 => x"842a8132",
  1190 => x"810657ff",
  1191 => x"537680f7",
  1192 => x"3873822a",
  1193 => x"70810651",
  1194 => x"5372802e",
  1195 => x"b938b015",
  1196 => x"08547380",
  1197 => x"2e9c3880",
  1198 => x"c0155373",
  1199 => x"732e8f38",
  1200 => x"735280cf",
  1201 => x"dc085187",
  1202 => x"ca3f8c15",
  1203 => x"225676b0",
  1204 => x"160c75db",
  1205 => x"0653728c",
  1206 => x"1623800b",
  1207 => x"84160c90",
  1208 => x"1508750c",
  1209 => x"72567588",
  1210 => x"0753728c",
  1211 => x"16239015",
  1212 => x"08802e80",
  1213 => x"c1388c15",
  1214 => x"22708106",
  1215 => x"5553739e",
  1216 => x"38720a10",
  1217 => x"0a708106",
  1218 => x"51537285",
  1219 => x"38941508",
  1220 => x"54738816",
  1221 => x"0c805372",
  1222 => x"800c883d",
  1223 => x"0d04800b",
  1224 => x"88160c94",
  1225 => x"15083098",
  1226 => x"160c8053",
  1227 => x"ea397251",
  1228 => x"82fb3ffe",
  1229 => x"c4397451",
  1230 => x"8ce83f8c",
  1231 => x"15227081",
  1232 => x"06555373",
  1233 => x"802effb9",
  1234 => x"38d439f8",
  1235 => x"3d0d7a58",
  1236 => x"77802e81",
  1237 => x"993880cf",
  1238 => x"dc0854b8",
  1239 => x"1408802e",
  1240 => x"80ed388c",
  1241 => x"18227090",
  1242 => x"2b70902c",
  1243 => x"70832a81",
  1244 => x"3281065c",
  1245 => x"51575478",
  1246 => x"80cd3890",
  1247 => x"18085776",
  1248 => x"802e80c3",
  1249 => x"38770877",
  1250 => x"3177790c",
  1251 => x"7683067a",
  1252 => x"58555573",
  1253 => x"85389418",
  1254 => x"08567588",
  1255 => x"190c8075",
  1256 => x"25a53874",
  1257 => x"5376529c",
  1258 => x"180851a4",
  1259 => x"18085473",
  1260 => x"2d800b80",
  1261 => x"082580c9",
  1262 => x"38800817",
  1263 => x"75800831",
  1264 => x"56577480",
  1265 => x"24dd3880",
  1266 => x"0b800c8a",
  1267 => x"3d0d0473",
  1268 => x"5181da3f",
  1269 => x"8c182270",
  1270 => x"902b7090",
  1271 => x"2c70832a",
  1272 => x"81328106",
  1273 => x"5c515754",
  1274 => x"78dd38ff",
  1275 => x"8e39a6cb",
  1276 => x"5280cfdc",
  1277 => x"085189f1",
  1278 => x"3f800880",
  1279 => x"0c8a3d0d",
  1280 => x"048c1822",
  1281 => x"80c00754",
  1282 => x"738c1923",
  1283 => x"ff0b800c",
  1284 => x"8a3d0d04",
  1285 => x"803d0d72",
  1286 => x"5180710c",
  1287 => x"800b8412",
  1288 => x"0c800b88",
  1289 => x"120c028e",
  1290 => x"05228c12",
  1291 => x"23029205",
  1292 => x"228e1223",
  1293 => x"800b9012",
  1294 => x"0c800b94",
  1295 => x"120c800b",
  1296 => x"98120c70",
  1297 => x"9c120c80",
  1298 => x"c2e00ba0",
  1299 => x"120c80c3",
  1300 => x"ac0ba412",
  1301 => x"0c80c4a8",
  1302 => x"0ba8120c",
  1303 => x"80c4f90b",
  1304 => x"ac120c82",
  1305 => x"3d0d04fa",
  1306 => x"3d0d7970",
  1307 => x"80dc298c",
  1308 => x"11547a53",
  1309 => x"56578cad",
  1310 => x"3f800880",
  1311 => x"08555680",
  1312 => x"08802ea2",
  1313 => x"3880088c",
  1314 => x"0554800b",
  1315 => x"80080c76",
  1316 => x"80088405",
  1317 => x"0c738008",
  1318 => x"88050c74",
  1319 => x"53805273",
  1320 => x"5197f83f",
  1321 => x"75547380",
  1322 => x"0c883d0d",
  1323 => x"04fc3d0d",
  1324 => x"76abc00b",
  1325 => x"bc120c55",
  1326 => x"810bb816",
  1327 => x"0c800b84",
  1328 => x"dc160c83",
  1329 => x"0b84e016",
  1330 => x"0c84e815",
  1331 => x"84e4160c",
  1332 => x"74548053",
  1333 => x"84528415",
  1334 => x"0851feb8",
  1335 => x"3f745481",
  1336 => x"53895288",
  1337 => x"150851fe",
  1338 => x"ab3f7454",
  1339 => x"82538a52",
  1340 => x"8c150851",
  1341 => x"fe9e3f86",
  1342 => x"3d0d04f9",
  1343 => x"3d0d7980",
  1344 => x"cfdc0854",
  1345 => x"57b81308",
  1346 => x"802e80c8",
  1347 => x"3884dc13",
  1348 => x"56881608",
  1349 => x"841708ff",
  1350 => x"05555580",
  1351 => x"74249f38",
  1352 => x"8c152270",
  1353 => x"902b7090",
  1354 => x"2c515458",
  1355 => x"72802e80",
  1356 => x"ca3880dc",
  1357 => x"15ff1555",
  1358 => x"55738025",
  1359 => x"e3387508",
  1360 => x"5372802e",
  1361 => x"9f387256",
  1362 => x"88160884",
  1363 => x"1708ff05",
  1364 => x"5555c839",
  1365 => x"7251fed5",
  1366 => x"3f80cfdc",
  1367 => x"0884dc05",
  1368 => x"56ffae39",
  1369 => x"84527651",
  1370 => x"fdfd3f80",
  1371 => x"08760c80",
  1372 => x"08802e80",
  1373 => x"c0388008",
  1374 => x"56ce3981",
  1375 => x"0b8c1623",
  1376 => x"72750c72",
  1377 => x"88160c72",
  1378 => x"84160c72",
  1379 => x"90160c72",
  1380 => x"94160c72",
  1381 => x"98160cff",
  1382 => x"0b8e1623",
  1383 => x"72b0160c",
  1384 => x"72b4160c",
  1385 => x"7280c416",
  1386 => x"0c7280c8",
  1387 => x"160c7480",
  1388 => x"0c893d0d",
  1389 => x"048c770c",
  1390 => x"800b800c",
  1391 => x"893d0d04",
  1392 => x"ff3d0da6",
  1393 => x"cb527351",
  1394 => x"869f3f83",
  1395 => x"3d0d0480",
  1396 => x"3d0d80cf",
  1397 => x"dc0851e8",
  1398 => x"3f823d0d",
  1399 => x"04fb3d0d",
  1400 => x"77705256",
  1401 => x"96c43f80",
  1402 => x"d7980b88",
  1403 => x"05088411",
  1404 => x"08fc0670",
  1405 => x"7b319fef",
  1406 => x"05e08006",
  1407 => x"e0800556",
  1408 => x"5653a080",
  1409 => x"74249438",
  1410 => x"80527551",
  1411 => x"969e3f80",
  1412 => x"d7a00815",
  1413 => x"53728008",
  1414 => x"2e8f3875",
  1415 => x"51968c3f",
  1416 => x"80537280",
  1417 => x"0c873d0d",
  1418 => x"04733052",
  1419 => x"755195fc",
  1420 => x"3f8008ff",
  1421 => x"2ea83880",
  1422 => x"d7980b88",
  1423 => x"05087575",
  1424 => x"31810784",
  1425 => x"120c5380",
  1426 => x"d6dc0874",
  1427 => x"3180d6dc",
  1428 => x"0c755195",
  1429 => x"d63f810b",
  1430 => x"800c873d",
  1431 => x"0d048052",
  1432 => x"755195c8",
  1433 => x"3f80d798",
  1434 => x"0b880508",
  1435 => x"80087131",
  1436 => x"56538f75",
  1437 => x"25ffa438",
  1438 => x"800880d7",
  1439 => x"8c083180",
  1440 => x"d6dc0c74",
  1441 => x"81078414",
  1442 => x"0c755195",
  1443 => x"9e3f8053",
  1444 => x"ff9039f6",
  1445 => x"3d0d7c7e",
  1446 => x"545b7280",
  1447 => x"2e828338",
  1448 => x"7a519586",
  1449 => x"3ff81384",
  1450 => x"110870fe",
  1451 => x"06701384",
  1452 => x"1108fc06",
  1453 => x"5d585954",
  1454 => x"5880d7a0",
  1455 => x"08752e82",
  1456 => x"de387884",
  1457 => x"160c8073",
  1458 => x"8106545a",
  1459 => x"727a2e81",
  1460 => x"d5387815",
  1461 => x"84110881",
  1462 => x"06515372",
  1463 => x"a0387817",
  1464 => x"577981e6",
  1465 => x"38881508",
  1466 => x"537280d7",
  1467 => x"a02e82f9",
  1468 => x"388c1508",
  1469 => x"708c150c",
  1470 => x"7388120c",
  1471 => x"56768107",
  1472 => x"84190c76",
  1473 => x"1877710c",
  1474 => x"53798191",
  1475 => x"3883ff77",
  1476 => x"2781c838",
  1477 => x"76892a77",
  1478 => x"832a5653",
  1479 => x"72802ebf",
  1480 => x"3876862a",
  1481 => x"b8055584",
  1482 => x"7327b438",
  1483 => x"80db1355",
  1484 => x"947327ab",
  1485 => x"38768c2a",
  1486 => x"80ee0555",
  1487 => x"80d47327",
  1488 => x"9e38768f",
  1489 => x"2a80f705",
  1490 => x"5582d473",
  1491 => x"27913876",
  1492 => x"922a80fc",
  1493 => x"05558ad4",
  1494 => x"73278438",
  1495 => x"80fe5574",
  1496 => x"10101080",
  1497 => x"d7980588",
  1498 => x"11085556",
  1499 => x"73762e82",
  1500 => x"b3388414",
  1501 => x"08fc0653",
  1502 => x"7673278d",
  1503 => x"38881408",
  1504 => x"5473762e",
  1505 => x"098106ea",
  1506 => x"388c1408",
  1507 => x"708c1a0c",
  1508 => x"74881a0c",
  1509 => x"7888120c",
  1510 => x"56778c15",
  1511 => x"0c7a5193",
  1512 => x"8a3f8c3d",
  1513 => x"0d047708",
  1514 => x"78713159",
  1515 => x"77058819",
  1516 => x"08545772",
  1517 => x"80d7a02e",
  1518 => x"80e0388c",
  1519 => x"1808708c",
  1520 => x"150c7388",
  1521 => x"120c56fe",
  1522 => x"89398815",
  1523 => x"088c1608",
  1524 => x"708c130c",
  1525 => x"5788170c",
  1526 => x"fea33976",
  1527 => x"832a7054",
  1528 => x"55807524",
  1529 => x"81983872",
  1530 => x"822c8171",
  1531 => x"2b80d79c",
  1532 => x"080780d7",
  1533 => x"980b8405",
  1534 => x"0c537410",
  1535 => x"101080d7",
  1536 => x"98058811",
  1537 => x"08555675",
  1538 => x"8c190c73",
  1539 => x"88190c77",
  1540 => x"88170c77",
  1541 => x"8c150cff",
  1542 => x"8439815a",
  1543 => x"fdb43978",
  1544 => x"17738106",
  1545 => x"54577298",
  1546 => x"38770878",
  1547 => x"71315977",
  1548 => x"058c1908",
  1549 => x"881a0871",
  1550 => x"8c120c88",
  1551 => x"120c5757",
  1552 => x"76810784",
  1553 => x"190c7780",
  1554 => x"d7980b88",
  1555 => x"050c80d7",
  1556 => x"94087726",
  1557 => x"fec73880",
  1558 => x"d7900852",
  1559 => x"7a51fafd",
  1560 => x"3f7a5191",
  1561 => x"c63ffeba",
  1562 => x"3981788c",
  1563 => x"150c7888",
  1564 => x"150c738c",
  1565 => x"1a0c7388",
  1566 => x"1a0c5afd",
  1567 => x"80398315",
  1568 => x"70822c81",
  1569 => x"712b80d7",
  1570 => x"9c080780",
  1571 => x"d7980b84",
  1572 => x"050c5153",
  1573 => x"74101010",
  1574 => x"80d79805",
  1575 => x"88110855",
  1576 => x"56fee439",
  1577 => x"74538075",
  1578 => x"24a73872",
  1579 => x"822c8171",
  1580 => x"2b80d79c",
  1581 => x"080780d7",
  1582 => x"980b8405",
  1583 => x"0c53758c",
  1584 => x"190c7388",
  1585 => x"190c7788",
  1586 => x"170c778c",
  1587 => x"150cfdcd",
  1588 => x"39831570",
  1589 => x"822c8171",
  1590 => x"2b80d79c",
  1591 => x"080780d7",
  1592 => x"980b8405",
  1593 => x"0c5153d6",
  1594 => x"39f93d0d",
  1595 => x"797b5853",
  1596 => x"800b80cf",
  1597 => x"dc085356",
  1598 => x"72722e80",
  1599 => x"c03884dc",
  1600 => x"13557476",
  1601 => x"2eb73888",
  1602 => x"15088416",
  1603 => x"08ff0554",
  1604 => x"54807324",
  1605 => x"9d388c14",
  1606 => x"2270902b",
  1607 => x"70902c51",
  1608 => x"53587180",
  1609 => x"d83880dc",
  1610 => x"14ff1454",
  1611 => x"54728025",
  1612 => x"e5387408",
  1613 => x"5574d038",
  1614 => x"80cfdc08",
  1615 => x"5284dc12",
  1616 => x"5574802e",
  1617 => x"b1388815",
  1618 => x"08841608",
  1619 => x"ff055454",
  1620 => x"8073249c",
  1621 => x"388c1422",
  1622 => x"70902b70",
  1623 => x"902c5153",
  1624 => x"5871ad38",
  1625 => x"80dc14ff",
  1626 => x"14545472",
  1627 => x"8025e638",
  1628 => x"74085574",
  1629 => x"d1387580",
  1630 => x"0c893d0d",
  1631 => x"04735176",
  1632 => x"2d758008",
  1633 => x"0780dc15",
  1634 => x"ff155555",
  1635 => x"56ff9e39",
  1636 => x"7351762d",
  1637 => x"75800807",
  1638 => x"80dc15ff",
  1639 => x"15555556",
  1640 => x"ca39ea3d",
  1641 => x"0d688c11",
  1642 => x"22700a10",
  1643 => x"0a810657",
  1644 => x"58567480",
  1645 => x"e4388e16",
  1646 => x"2270902b",
  1647 => x"70902c51",
  1648 => x"55588074",
  1649 => x"24b13898",
  1650 => x"3dc40553",
  1651 => x"735280cf",
  1652 => x"dc085192",
  1653 => x"ac3f800b",
  1654 => x"80082497",
  1655 => x"387983e0",
  1656 => x"80065473",
  1657 => x"80c0802e",
  1658 => x"818f3873",
  1659 => x"8280802e",
  1660 => x"8191388c",
  1661 => x"16225776",
  1662 => x"90800754",
  1663 => x"738c1723",
  1664 => x"88805280",
  1665 => x"cfdc0851",
  1666 => x"819b3f80",
  1667 => x"089d388c",
  1668 => x"16228207",
  1669 => x"54738c17",
  1670 => x"2380c316",
  1671 => x"70770c90",
  1672 => x"170c810b",
  1673 => x"94170c98",
  1674 => x"3d0d0480",
  1675 => x"cfdc08ab",
  1676 => x"c00bbc12",
  1677 => x"0c548c16",
  1678 => x"22818007",
  1679 => x"54738c17",
  1680 => x"23800876",
  1681 => x"0c800890",
  1682 => x"170c8880",
  1683 => x"0b94170c",
  1684 => x"74802ed3",
  1685 => x"388e1622",
  1686 => x"70902b70",
  1687 => x"902c5355",
  1688 => x"5898aa3f",
  1689 => x"8008802e",
  1690 => x"ffbd388c",
  1691 => x"16228107",
  1692 => x"54738c17",
  1693 => x"23983d0d",
  1694 => x"04810b8c",
  1695 => x"17225855",
  1696 => x"fef539a8",
  1697 => x"160880c4",
  1698 => x"a82e0981",
  1699 => x"06fee438",
  1700 => x"8c162288",
  1701 => x"80075473",
  1702 => x"8c172388",
  1703 => x"800b80cc",
  1704 => x"170cfedc",
  1705 => x"39f33d0d",
  1706 => x"7f618b11",
  1707 => x"70f8065c",
  1708 => x"55555e72",
  1709 => x"96268338",
  1710 => x"90598079",
  1711 => x"24747a26",
  1712 => x"07538054",
  1713 => x"72742e09",
  1714 => x"810680cb",
  1715 => x"387d518c",
  1716 => x"d93f7883",
  1717 => x"f72680c6",
  1718 => x"3878832a",
  1719 => x"70101010",
  1720 => x"80d79805",
  1721 => x"8c110859",
  1722 => x"595a7678",
  1723 => x"2e83b038",
  1724 => x"841708fc",
  1725 => x"06568c17",
  1726 => x"08881808",
  1727 => x"718c120c",
  1728 => x"88120c58",
  1729 => x"75178411",
  1730 => x"08810784",
  1731 => x"120c537d",
  1732 => x"518c983f",
  1733 => x"88175473",
  1734 => x"800c8f3d",
  1735 => x"0d047889",
  1736 => x"2a79832a",
  1737 => x"5b537280",
  1738 => x"2ebf3878",
  1739 => x"862ab805",
  1740 => x"5a847327",
  1741 => x"b43880db",
  1742 => x"135a9473",
  1743 => x"27ab3878",
  1744 => x"8c2a80ee",
  1745 => x"055a80d4",
  1746 => x"73279e38",
  1747 => x"788f2a80",
  1748 => x"f7055a82",
  1749 => x"d4732791",
  1750 => x"3878922a",
  1751 => x"80fc055a",
  1752 => x"8ad47327",
  1753 => x"843880fe",
  1754 => x"5a791010",
  1755 => x"1080d798",
  1756 => x"058c1108",
  1757 => x"58557675",
  1758 => x"2ea33884",
  1759 => x"1708fc06",
  1760 => x"707a3155",
  1761 => x"56738f24",
  1762 => x"88d53873",
  1763 => x"8025fee6",
  1764 => x"388c1708",
  1765 => x"5776752e",
  1766 => x"098106df",
  1767 => x"38811a5a",
  1768 => x"80d7a808",
  1769 => x"577680d7",
  1770 => x"a02e82c0",
  1771 => x"38841708",
  1772 => x"fc06707a",
  1773 => x"31555673",
  1774 => x"8f2481f9",
  1775 => x"3880d7a0",
  1776 => x"0b80d7ac",
  1777 => x"0c80d7a0",
  1778 => x"0b80d7a8",
  1779 => x"0c738025",
  1780 => x"feb23883",
  1781 => x"ff762783",
  1782 => x"df387589",
  1783 => x"2a76832a",
  1784 => x"55537280",
  1785 => x"2ebf3875",
  1786 => x"862ab805",
  1787 => x"54847327",
  1788 => x"b43880db",
  1789 => x"13549473",
  1790 => x"27ab3875",
  1791 => x"8c2a80ee",
  1792 => x"055480d4",
  1793 => x"73279e38",
  1794 => x"758f2a80",
  1795 => x"f7055482",
  1796 => x"d4732791",
  1797 => x"3875922a",
  1798 => x"80fc0554",
  1799 => x"8ad47327",
  1800 => x"843880fe",
  1801 => x"54731010",
  1802 => x"1080d798",
  1803 => x"05881108",
  1804 => x"56587478",
  1805 => x"2e86cf38",
  1806 => x"841508fc",
  1807 => x"06537573",
  1808 => x"278d3888",
  1809 => x"15085574",
  1810 => x"782e0981",
  1811 => x"06ea388c",
  1812 => x"150880d7",
  1813 => x"980b8405",
  1814 => x"08718c1a",
  1815 => x"0c76881a",
  1816 => x"0c788813",
  1817 => x"0c788c18",
  1818 => x"0c5d5879",
  1819 => x"53807a24",
  1820 => x"83e63872",
  1821 => x"822c8171",
  1822 => x"2b5c537a",
  1823 => x"7c268198",
  1824 => x"387b7b06",
  1825 => x"537282f1",
  1826 => x"3879fc06",
  1827 => x"84055a7a",
  1828 => x"10707d06",
  1829 => x"545b7282",
  1830 => x"e038841a",
  1831 => x"5af13988",
  1832 => x"178c1108",
  1833 => x"58587678",
  1834 => x"2e098106",
  1835 => x"fcc23882",
  1836 => x"1a5afdec",
  1837 => x"39781779",
  1838 => x"81078419",
  1839 => x"0c7080d7",
  1840 => x"ac0c7080",
  1841 => x"d7a80c80",
  1842 => x"d7a00b8c",
  1843 => x"120c8c11",
  1844 => x"0888120c",
  1845 => x"74810784",
  1846 => x"120c7411",
  1847 => x"75710c51",
  1848 => x"537d5188",
  1849 => x"c63f8817",
  1850 => x"54fcac39",
  1851 => x"80d7980b",
  1852 => x"8405087a",
  1853 => x"545c7980",
  1854 => x"25fef838",
  1855 => x"82da397a",
  1856 => x"097c0670",
  1857 => x"80d7980b",
  1858 => x"84050c5c",
  1859 => x"7a105b7a",
  1860 => x"7c268538",
  1861 => x"7a85b838",
  1862 => x"80d7980b",
  1863 => x"88050870",
  1864 => x"841208fc",
  1865 => x"06707c31",
  1866 => x"7c72268f",
  1867 => x"72250757",
  1868 => x"575c5d55",
  1869 => x"72802e80",
  1870 => x"db38797a",
  1871 => x"1680d790",
  1872 => x"081b9011",
  1873 => x"5a55575b",
  1874 => x"80d78c08",
  1875 => x"ff2e8838",
  1876 => x"a08f13e0",
  1877 => x"80065776",
  1878 => x"527d5187",
  1879 => x"cf3f8008",
  1880 => x"548008ff",
  1881 => x"2e903880",
  1882 => x"08762782",
  1883 => x"99387480",
  1884 => x"d7982e82",
  1885 => x"913880d7",
  1886 => x"980b8805",
  1887 => x"08558415",
  1888 => x"08fc0670",
  1889 => x"7a317a72",
  1890 => x"268f7225",
  1891 => x"07525553",
  1892 => x"7283e638",
  1893 => x"74798107",
  1894 => x"84170c79",
  1895 => x"167080d7",
  1896 => x"980b8805",
  1897 => x"0c758107",
  1898 => x"84120c54",
  1899 => x"7e525786",
  1900 => x"fa3f8817",
  1901 => x"54fae039",
  1902 => x"75832a70",
  1903 => x"54548074",
  1904 => x"24819b38",
  1905 => x"72822c81",
  1906 => x"712b80d7",
  1907 => x"9c080770",
  1908 => x"80d7980b",
  1909 => x"84050c75",
  1910 => x"10101080",
  1911 => x"d7980588",
  1912 => x"1108585a",
  1913 => x"5d53778c",
  1914 => x"180c7488",
  1915 => x"180c7688",
  1916 => x"190c768c",
  1917 => x"160cfcf3",
  1918 => x"39797a10",
  1919 => x"101080d7",
  1920 => x"98057057",
  1921 => x"595d8c15",
  1922 => x"08577675",
  1923 => x"2ea33884",
  1924 => x"1708fc06",
  1925 => x"707a3155",
  1926 => x"56738f24",
  1927 => x"83ca3873",
  1928 => x"80258481",
  1929 => x"388c1708",
  1930 => x"5776752e",
  1931 => x"098106df",
  1932 => x"38881581",
  1933 => x"1b708306",
  1934 => x"555b5572",
  1935 => x"c9387c83",
  1936 => x"06537280",
  1937 => x"2efdb838",
  1938 => x"ff1df819",
  1939 => x"595d8818",
  1940 => x"08782eea",
  1941 => x"38fdb539",
  1942 => x"831a53fc",
  1943 => x"96398314",
  1944 => x"70822c81",
  1945 => x"712b80d7",
  1946 => x"9c080770",
  1947 => x"80d7980b",
  1948 => x"84050c76",
  1949 => x"10101080",
  1950 => x"d7980588",
  1951 => x"1108595b",
  1952 => x"5e5153fe",
  1953 => x"e13980d6",
  1954 => x"dc081758",
  1955 => x"8008762e",
  1956 => x"818d3880",
  1957 => x"d78c08ff",
  1958 => x"2e83ec38",
  1959 => x"73763118",
  1960 => x"80d6dc0c",
  1961 => x"73870670",
  1962 => x"57537280",
  1963 => x"2e883888",
  1964 => x"73317015",
  1965 => x"55567614",
  1966 => x"9fff06a0",
  1967 => x"80713117",
  1968 => x"70547f53",
  1969 => x"575384e4",
  1970 => x"3f800853",
  1971 => x"8008ff2e",
  1972 => x"81a03880",
  1973 => x"d6dc0816",
  1974 => x"7080d6dc",
  1975 => x"0c747580",
  1976 => x"d7980b88",
  1977 => x"050c7476",
  1978 => x"31187081",
  1979 => x"07515556",
  1980 => x"587b80d7",
  1981 => x"982e839c",
  1982 => x"38798f26",
  1983 => x"82cb3881",
  1984 => x"0b84150c",
  1985 => x"841508fc",
  1986 => x"06707a31",
  1987 => x"7a72268f",
  1988 => x"72250752",
  1989 => x"55537280",
  1990 => x"2efcf938",
  1991 => x"80db3980",
  1992 => x"089fff06",
  1993 => x"5372feeb",
  1994 => x"387780d6",
  1995 => x"dc0c80d7",
  1996 => x"980b8805",
  1997 => x"087b1881",
  1998 => x"0784120c",
  1999 => x"5580d788",
  2000 => x"08782786",
  2001 => x"387780d7",
  2002 => x"880c80d7",
  2003 => x"84087827",
  2004 => x"fcac3877",
  2005 => x"80d7840c",
  2006 => x"841508fc",
  2007 => x"06707a31",
  2008 => x"7a72268f",
  2009 => x"72250752",
  2010 => x"55537280",
  2011 => x"2efca538",
  2012 => x"88398074",
  2013 => x"5456fedb",
  2014 => x"397d5183",
  2015 => x"ae3f800b",
  2016 => x"800c8f3d",
  2017 => x"0d047353",
  2018 => x"807424a9",
  2019 => x"3872822c",
  2020 => x"81712b80",
  2021 => x"d79c0807",
  2022 => x"7080d798",
  2023 => x"0b84050c",
  2024 => x"5d53778c",
  2025 => x"180c7488",
  2026 => x"180c7688",
  2027 => x"190c768c",
  2028 => x"160cf9b7",
  2029 => x"39831470",
  2030 => x"822c8171",
  2031 => x"2b80d79c",
  2032 => x"08077080",
  2033 => x"d7980b84",
  2034 => x"050c5e51",
  2035 => x"53d4397b",
  2036 => x"7b065372",
  2037 => x"fca33884",
  2038 => x"1a7b105c",
  2039 => x"5af139ff",
  2040 => x"1a811151",
  2041 => x"5af7b939",
  2042 => x"78177981",
  2043 => x"0784190c",
  2044 => x"8c180888",
  2045 => x"1908718c",
  2046 => x"120c8812",
  2047 => x"0c597080",
  2048 => x"d7ac0c70",
  2049 => x"80d7a80c",
  2050 => x"80d7a00b",
  2051 => x"8c120c8c",
  2052 => x"11088812",
  2053 => x"0c748107",
  2054 => x"84120c74",
  2055 => x"1175710c",
  2056 => x"5153f9bd",
  2057 => x"39751784",
  2058 => x"11088107",
  2059 => x"84120c53",
  2060 => x"8c170888",
  2061 => x"1808718c",
  2062 => x"120c8812",
  2063 => x"0c587d51",
  2064 => x"81e93f88",
  2065 => x"1754f5cf",
  2066 => x"39728415",
  2067 => x"0cf41af8",
  2068 => x"0670841e",
  2069 => x"08810607",
  2070 => x"841e0c70",
  2071 => x"1d545b85",
  2072 => x"0b84140c",
  2073 => x"850b8814",
  2074 => x"0c8f7b27",
  2075 => x"fdcf3888",
  2076 => x"1c527d51",
  2077 => x"ec9d3f80",
  2078 => x"d7980b88",
  2079 => x"050880d6",
  2080 => x"dc085955",
  2081 => x"fdb73977",
  2082 => x"80d6dc0c",
  2083 => x"7380d78c",
  2084 => x"0cfc9139",
  2085 => x"7284150c",
  2086 => x"fda339fc",
  2087 => x"3d0d7679",
  2088 => x"71028c05",
  2089 => x"9f053357",
  2090 => x"55535583",
  2091 => x"72278a38",
  2092 => x"74830651",
  2093 => x"70802ea2",
  2094 => x"38ff1252",
  2095 => x"71ff2e93",
  2096 => x"38737370",
  2097 => x"81055534",
  2098 => x"ff125271",
  2099 => x"ff2e0981",
  2100 => x"06ef3874",
  2101 => x"800c863d",
  2102 => x"0d047474",
  2103 => x"882b7507",
  2104 => x"7071902b",
  2105 => x"07515451",
  2106 => x"8f7227a5",
  2107 => x"38727170",
  2108 => x"8405530c",
  2109 => x"72717084",
  2110 => x"05530c72",
  2111 => x"71708405",
  2112 => x"530c7271",
  2113 => x"70840553",
  2114 => x"0cf01252",
  2115 => x"718f26dd",
  2116 => x"38837227",
  2117 => x"90387271",
  2118 => x"70840553",
  2119 => x"0cfc1252",
  2120 => x"718326f2",
  2121 => x"387053ff",
  2122 => x"90390404",
  2123 => x"fd3d0d80",
  2124 => x"0b80dfd0",
  2125 => x"0c765184",
  2126 => x"ee3f8008",
  2127 => x"538008ff",
  2128 => x"2e883872",
  2129 => x"800c853d",
  2130 => x"0d0480df",
  2131 => x"d0085473",
  2132 => x"802ef038",
  2133 => x"7574710c",
  2134 => x"5272800c",
  2135 => x"853d0d04",
  2136 => x"f93d0d79",
  2137 => x"7c557b54",
  2138 => x"8e112270",
  2139 => x"902b7090",
  2140 => x"2c555780",
  2141 => x"cfdc0853",
  2142 => x"585683f3",
  2143 => x"3f800857",
  2144 => x"800b8008",
  2145 => x"24933880",
  2146 => x"d0160880",
  2147 => x"080580d0",
  2148 => x"170c7680",
  2149 => x"0c893d0d",
  2150 => x"048c1622",
  2151 => x"83dfff06",
  2152 => x"55748c17",
  2153 => x"2376800c",
  2154 => x"893d0d04",
  2155 => x"fa3d0d78",
  2156 => x"8c112270",
  2157 => x"882a7081",
  2158 => x"06515758",
  2159 => x"5674a938",
  2160 => x"8c162283",
  2161 => x"dfff0655",
  2162 => x"748c1723",
  2163 => x"7a547953",
  2164 => x"8e162270",
  2165 => x"902b7090",
  2166 => x"2c545680",
  2167 => x"cfdc0852",
  2168 => x"5681b23f",
  2169 => x"883d0d04",
  2170 => x"82548053",
  2171 => x"8e162270",
  2172 => x"902b7090",
  2173 => x"2c545680",
  2174 => x"cfdc0852",
  2175 => x"5782b83f",
  2176 => x"8c162283",
  2177 => x"dfff0655",
  2178 => x"748c1723",
  2179 => x"7a547953",
  2180 => x"8e162270",
  2181 => x"902b7090",
  2182 => x"2c545680",
  2183 => x"cfdc0852",
  2184 => x"5680f23f",
  2185 => x"883d0d04",
  2186 => x"f93d0d79",
  2187 => x"7c557b54",
  2188 => x"8e112270",
  2189 => x"902b7090",
  2190 => x"2c555780",
  2191 => x"cfdc0853",
  2192 => x"585681f3",
  2193 => x"3f800857",
  2194 => x"8008ff2e",
  2195 => x"99388c16",
  2196 => x"22a08007",
  2197 => x"55748c17",
  2198 => x"23800880",
  2199 => x"d0170c76",
  2200 => x"800c893d",
  2201 => x"0d048c16",
  2202 => x"2283dfff",
  2203 => x"0655748c",
  2204 => x"17237680",
  2205 => x"0c893d0d",
  2206 => x"04fe3d0d",
  2207 => x"748e1122",
  2208 => x"70902b70",
  2209 => x"902c5551",
  2210 => x"515380cf",
  2211 => x"dc0851bd",
  2212 => x"3f843d0d",
  2213 => x"04fb3d0d",
  2214 => x"800b80df",
  2215 => x"d00c7a53",
  2216 => x"79527851",
  2217 => x"82fd3f80",
  2218 => x"08558008",
  2219 => x"ff2e8838",
  2220 => x"74800c87",
  2221 => x"3d0d0480",
  2222 => x"dfd00856",
  2223 => x"75802ef0",
  2224 => x"38777671",
  2225 => x"0c547480",
  2226 => x"0c873d0d",
  2227 => x"04fd3d0d",
  2228 => x"800b80df",
  2229 => x"d00c7651",
  2230 => x"84cc3f80",
  2231 => x"08538008",
  2232 => x"ff2e8838",
  2233 => x"72800c85",
  2234 => x"3d0d0480",
  2235 => x"dfd00854",
  2236 => x"73802ef0",
  2237 => x"38757471",
  2238 => x"0c527280",
  2239 => x"0c853d0d",
  2240 => x"04fc3d0d",
  2241 => x"800b80df",
  2242 => x"d00c7852",
  2243 => x"775186b4",
  2244 => x"3f800854",
  2245 => x"8008ff2e",
  2246 => x"88387380",
  2247 => x"0c863d0d",
  2248 => x"0480dfd0",
  2249 => x"08557480",
  2250 => x"2ef03876",
  2251 => x"75710c53",
  2252 => x"73800c86",
  2253 => x"3d0d04fb",
  2254 => x"3d0d800b",
  2255 => x"80dfd00c",
  2256 => x"7a537952",
  2257 => x"78518490",
  2258 => x"3f800855",
  2259 => x"8008ff2e",
  2260 => x"88387480",
  2261 => x"0c873d0d",
  2262 => x"0480dfd0",
  2263 => x"08567580",
  2264 => x"2ef03877",
  2265 => x"76710c54",
  2266 => x"74800c87",
  2267 => x"3d0d04fb",
  2268 => x"3d0d800b",
  2269 => x"80dfd00c",
  2270 => x"7a537952",
  2271 => x"78518298",
  2272 => x"3f800855",
  2273 => x"8008ff2e",
  2274 => x"88387480",
  2275 => x"0c873d0d",
  2276 => x"0480dfd0",
  2277 => x"08567580",
  2278 => x"2ef03877",
  2279 => x"76710c54",
  2280 => x"74800c87",
  2281 => x"3d0d04fe",
  2282 => x"3d0d80df",
  2283 => x"c8085170",
  2284 => x"8a3880df",
  2285 => x"d47080df",
  2286 => x"c80c5170",
  2287 => x"75125252",
  2288 => x"ff537087",
  2289 => x"fb808026",
  2290 => x"88387080",
  2291 => x"dfc80c71",
  2292 => x"5372800c",
  2293 => x"843d0d04",
  2294 => x"fd3d0d80",
  2295 => x"0b80cfd0",
  2296 => x"08545472",
  2297 => x"812e9b38",
  2298 => x"7380dfcc",
  2299 => x"0cc2ab3f",
  2300 => x"c08e3f80",
  2301 => x"dfa05281",
  2302 => x"51c1ca3f",
  2303 => x"80085185",
  2304 => x"c33f7280",
  2305 => x"dfcc0cc2",
  2306 => x"913fffbf",
  2307 => x"f33f80df",
  2308 => x"a0528151",
  2309 => x"c1af3f80",
  2310 => x"085185a8",
  2311 => x"3f00ff39",
  2312 => x"00ff39f5",
  2313 => x"3d0d7e60",
  2314 => x"80dfcc08",
  2315 => x"705b585b",
  2316 => x"5b7580c2",
  2317 => x"38777a25",
  2318 => x"a138771b",
  2319 => x"70337081",
  2320 => x"ff065858",
  2321 => x"59758a2e",
  2322 => x"98387681",
  2323 => x"ff0651c1",
  2324 => x"aa3f8118",
  2325 => x"58797824",
  2326 => x"e1387980",
  2327 => x"0c8d3d0d",
  2328 => x"048d51c1",
  2329 => x"963f7833",
  2330 => x"7081ff06",
  2331 => x"5257c18b",
  2332 => x"3f811858",
  2333 => x"e0397955",
  2334 => x"7a547d53",
  2335 => x"85528d3d",
  2336 => x"fc0551ff",
  2337 => x"bfbc3f80",
  2338 => x"085684b1",
  2339 => x"3f7b8008",
  2340 => x"0c75800c",
  2341 => x"8d3d0d04",
  2342 => x"f63d0d7d",
  2343 => x"7f80dfcc",
  2344 => x"08705b58",
  2345 => x"5a5a7580",
  2346 => x"c1387779",
  2347 => x"25b338c0",
  2348 => x"a73f8008",
  2349 => x"81ff0670",
  2350 => x"8d327030",
  2351 => x"709f2a51",
  2352 => x"51575776",
  2353 => x"8a2e80c4",
  2354 => x"3875802e",
  2355 => x"bf38771a",
  2356 => x"56767634",
  2357 => x"7651c0a3",
  2358 => x"3f811858",
  2359 => x"787824cf",
  2360 => x"38775675",
  2361 => x"800c8c3d",
  2362 => x"0d047855",
  2363 => x"79547c53",
  2364 => x"84528c3d",
  2365 => x"fc0551ff",
  2366 => x"bec83f80",
  2367 => x"085683bd",
  2368 => x"3f7a8008",
  2369 => x"0c75800c",
  2370 => x"8c3d0d04",
  2371 => x"771a568a",
  2372 => x"76348118",
  2373 => x"588d51ff",
  2374 => x"bfe13f8a",
  2375 => x"51ffbfdb",
  2376 => x"3f7756ff",
  2377 => x"be39fb3d",
  2378 => x"0d80dfcc",
  2379 => x"08705654",
  2380 => x"73883874",
  2381 => x"800c873d",
  2382 => x"0d047753",
  2383 => x"8352873d",
  2384 => x"fc0551ff",
  2385 => x"bdfc3f80",
  2386 => x"085482f1",
  2387 => x"3f758008",
  2388 => x"0c73800c",
  2389 => x"873d0d04",
  2390 => x"fa3d0d80",
  2391 => x"dfcc0880",
  2392 => x"2ea3387a",
  2393 => x"55795478",
  2394 => x"53865288",
  2395 => x"3dfc0551",
  2396 => x"ffbdcf3f",
  2397 => x"80085682",
  2398 => x"c43f7680",
  2399 => x"080c7580",
  2400 => x"0c883d0d",
  2401 => x"0482b63f",
  2402 => x"9d0b8008",
  2403 => x"0cff0b80",
  2404 => x"0c883d0d",
  2405 => x"04fb3d0d",
  2406 => x"77795656",
  2407 => x"80705454",
  2408 => x"7375259f",
  2409 => x"38741010",
  2410 => x"10f80552",
  2411 => x"72167033",
  2412 => x"70742b76",
  2413 => x"078116f8",
  2414 => x"16565656",
  2415 => x"51517473",
  2416 => x"24ea3873",
  2417 => x"800c873d",
  2418 => x"0d04fc3d",
  2419 => x"0d767855",
  2420 => x"55bc5380",
  2421 => x"527351f5",
  2422 => x"c23f8452",
  2423 => x"7451ffb5",
  2424 => x"3f800874",
  2425 => x"23845284",
  2426 => x"1551ffa9",
  2427 => x"3f800882",
  2428 => x"15238452",
  2429 => x"881551ff",
  2430 => x"9c3f8008",
  2431 => x"84150c84",
  2432 => x"528c1551",
  2433 => x"ff8f3f80",
  2434 => x"08881523",
  2435 => x"84529015",
  2436 => x"51ff823f",
  2437 => x"80088a15",
  2438 => x"23845294",
  2439 => x"1551fef5",
  2440 => x"3f80088c",
  2441 => x"15238452",
  2442 => x"981551fe",
  2443 => x"e83f8008",
  2444 => x"8e152388",
  2445 => x"529c1551",
  2446 => x"fedb3f80",
  2447 => x"0890150c",
  2448 => x"863d0d04",
  2449 => x"e93d0d6a",
  2450 => x"80dfcc08",
  2451 => x"57577593",
  2452 => x"3880c080",
  2453 => x"0b84180c",
  2454 => x"75ac180c",
  2455 => x"75800c99",
  2456 => x"3d0d0489",
  2457 => x"3d70556a",
  2458 => x"54558a52",
  2459 => x"993dffbc",
  2460 => x"0551ffbb",
  2461 => x"cd3f8008",
  2462 => x"77537552",
  2463 => x"56fecb3f",
  2464 => x"bc3f7780",
  2465 => x"080c7580",
  2466 => x"0c993d0d",
  2467 => x"04fc3d0d",
  2468 => x"815480df",
  2469 => x"cc088838",
  2470 => x"73800c86",
  2471 => x"3d0d0476",
  2472 => x"5397b952",
  2473 => x"863dfc05",
  2474 => x"51ffbb96",
  2475 => x"3f800854",
  2476 => x"8c3f7480",
  2477 => x"080c7380",
  2478 => x"0c863d0d",
  2479 => x"0480cfdc",
  2480 => x"08800c04",
  2481 => x"f73d0d7b",
  2482 => x"80cfdc08",
  2483 => x"82c81108",
  2484 => x"5a545a77",
  2485 => x"802e80da",
  2486 => x"38818818",
  2487 => x"841908ff",
  2488 => x"0581712b",
  2489 => x"59555980",
  2490 => x"742480ea",
  2491 => x"38807424",
  2492 => x"b5387382",
  2493 => x"2b781188",
  2494 => x"05565681",
  2495 => x"80190877",
  2496 => x"06537280",
  2497 => x"2eb63878",
  2498 => x"16700853",
  2499 => x"53795174",
  2500 => x"0853722d",
  2501 => x"ff14fc17",
  2502 => x"fc177981",
  2503 => x"2c5a5757",
  2504 => x"54738025",
  2505 => x"d6387708",
  2506 => x"5877ffad",
  2507 => x"3880cfdc",
  2508 => x"0853bc13",
  2509 => x"08a53879",
  2510 => x"51f9e23f",
  2511 => x"74085372",
  2512 => x"2dff14fc",
  2513 => x"17fc1779",
  2514 => x"812c5a57",
  2515 => x"57547380",
  2516 => x"25ffa838",
  2517 => x"d1398057",
  2518 => x"ff933972",
  2519 => x"51bc1308",
  2520 => x"53722d79",
  2521 => x"51f9b63f",
  2522 => x"ff3d0d80",
  2523 => x"dfa80bfc",
  2524 => x"05700852",
  2525 => x"5270ff2e",
  2526 => x"9138702d",
  2527 => x"fc127008",
  2528 => x"525270ff",
  2529 => x"2e098106",
  2530 => x"f138833d",
  2531 => x"0d0404ff",
  2532 => x"b9ce3f04",
  2533 => x"48656c6c",
  2534 => x"6f20776f",
  2535 => x"726c6421",
  2536 => x"00000000",
  2537 => x"00000040",
  2538 => x"0a000000",
  2539 => x"43000000",
  2540 => x"64756d6d",
  2541 => x"792e6578",
  2542 => x"65000000",
  2543 => x"00ffffff",
  2544 => x"ff00ffff",
  2545 => x"ffff00ff",
  2546 => x"ffffff00",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000000",
  2550 => x"00002fb0",
  2551 => x"000027e0",
  2552 => x"00000000",
  2553 => x"00002a48",
  2554 => x"00002aa4",
  2555 => x"00002b00",
  2556 => x"00000000",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"00000000",
  2560 => x"00000000",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000000",
  2564 => x"00000000",
  2565 => x"000027ac",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"00000000",
  2569 => x"00000000",
  2570 => x"00000000",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"00000000",
  2574 => x"00000000",
  2575 => x"00000000",
  2576 => x"00000000",
  2577 => x"00000000",
  2578 => x"00000000",
  2579 => x"00000000",
  2580 => x"00000000",
  2581 => x"00000000",
  2582 => x"00000000",
  2583 => x"00000000",
  2584 => x"00000000",
  2585 => x"00000000",
  2586 => x"00000000",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000000",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000000",
  2594 => x"00000001",
  2595 => x"330eabcd",
  2596 => x"1234e66d",
  2597 => x"deec0005",
  2598 => x"000b0000",
  2599 => x"00000000",
  2600 => x"00000000",
  2601 => x"00000000",
  2602 => x"00000000",
  2603 => x"00000000",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00000000",
  2607 => x"00000000",
  2608 => x"00000000",
  2609 => x"00000000",
  2610 => x"00000000",
  2611 => x"00000000",
  2612 => x"00000000",
  2613 => x"00000000",
  2614 => x"00000000",
  2615 => x"00000000",
  2616 => x"00000000",
  2617 => x"00000000",
  2618 => x"00000000",
  2619 => x"00000000",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000000",
  2623 => x"00000000",
  2624 => x"00000000",
  2625 => x"00000000",
  2626 => x"00000000",
  2627 => x"00000000",
  2628 => x"00000000",
  2629 => x"00000000",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000000",
  2633 => x"00000000",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00000000",
  2638 => x"00000000",
  2639 => x"00000000",
  2640 => x"00000000",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"00000000",
  2645 => x"00000000",
  2646 => x"00000000",
  2647 => x"00000000",
  2648 => x"00000000",
  2649 => x"00000000",
  2650 => x"00000000",
  2651 => x"00000000",
  2652 => x"00000000",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000000",
  2659 => x"00000000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"00000000",
  2715 => x"00000000",
  2716 => x"00000000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"00000000",
  2720 => x"00000000",
  2721 => x"00000000",
  2722 => x"00000000",
  2723 => x"00000000",
  2724 => x"00000000",
  2725 => x"00000000",
  2726 => x"00000000",
  2727 => x"00000000",
  2728 => x"00000000",
  2729 => x"00000000",
  2730 => x"00000000",
  2731 => x"00000000",
  2732 => x"00000000",
  2733 => x"00000000",
  2734 => x"00000000",
  2735 => x"00000000",
  2736 => x"00000000",
  2737 => x"00000000",
  2738 => x"00000000",
  2739 => x"00000000",
  2740 => x"00000000",
  2741 => x"00000000",
  2742 => x"00000000",
  2743 => x"00000000",
  2744 => x"00000000",
  2745 => x"00000000",
  2746 => x"00000000",
  2747 => x"00000000",
  2748 => x"00000000",
  2749 => x"00000000",
  2750 => x"00000000",
  2751 => x"00000000",
  2752 => x"00000000",
  2753 => x"00000000",
  2754 => x"00000000",
  2755 => x"00000000",
  2756 => x"00000000",
  2757 => x"00000000",
  2758 => x"00000000",
  2759 => x"00000000",
  2760 => x"00000000",
  2761 => x"00000000",
  2762 => x"00000000",
  2763 => x"00000000",
  2764 => x"00000000",
  2765 => x"00000000",
  2766 => x"00000000",
  2767 => x"00000000",
  2768 => x"00000000",
  2769 => x"00000000",
  2770 => x"00000000",
  2771 => x"00000000",
  2772 => x"00000000",
  2773 => x"00000000",
  2774 => x"00000000",
  2775 => x"00000000",
  2776 => x"00000000",
  2777 => x"00000000",
  2778 => x"00000000",
  2779 => x"00000000",
  2780 => x"00000000",
  2781 => x"00000000",
  2782 => x"00000000",
  2783 => x"00000000",
  2784 => x"00000000",
  2785 => x"00000000",
  2786 => x"00000000",
  2787 => x"ffffffff",
  2788 => x"00000000",
  2789 => x"00020000",
  2790 => x"00000000",
  2791 => x"00000000",
  2792 => x"00002b98",
  2793 => x"00002b98",
  2794 => x"00002ba0",
  2795 => x"00002ba0",
  2796 => x"00002ba8",
  2797 => x"00002ba8",
  2798 => x"00002bb0",
  2799 => x"00002bb0",
  2800 => x"00002bb8",
  2801 => x"00002bb8",
  2802 => x"00002bc0",
  2803 => x"00002bc0",
  2804 => x"00002bc8",
  2805 => x"00002bc8",
  2806 => x"00002bd0",
  2807 => x"00002bd0",
  2808 => x"00002bd8",
  2809 => x"00002bd8",
  2810 => x"00002be0",
  2811 => x"00002be0",
  2812 => x"00002be8",
  2813 => x"00002be8",
  2814 => x"00002bf0",
  2815 => x"00002bf0",
  2816 => x"00002bf8",
  2817 => x"00002bf8",
  2818 => x"00002c00",
  2819 => x"00002c00",
  2820 => x"00002c08",
  2821 => x"00002c08",
  2822 => x"00002c10",
  2823 => x"00002c10",
  2824 => x"00002c18",
  2825 => x"00002c18",
  2826 => x"00002c20",
  2827 => x"00002c20",
  2828 => x"00002c28",
  2829 => x"00002c28",
  2830 => x"00002c30",
  2831 => x"00002c30",
  2832 => x"00002c38",
  2833 => x"00002c38",
  2834 => x"00002c40",
  2835 => x"00002c40",
  2836 => x"00002c48",
  2837 => x"00002c48",
  2838 => x"00002c50",
  2839 => x"00002c50",
  2840 => x"00002c58",
  2841 => x"00002c58",
  2842 => x"00002c60",
  2843 => x"00002c60",
  2844 => x"00002c68",
  2845 => x"00002c68",
  2846 => x"00002c70",
  2847 => x"00002c70",
  2848 => x"00002c78",
  2849 => x"00002c78",
  2850 => x"00002c80",
  2851 => x"00002c80",
  2852 => x"00002c88",
  2853 => x"00002c88",
  2854 => x"00002c90",
  2855 => x"00002c90",
  2856 => x"00002c98",
  2857 => x"00002c98",
  2858 => x"00002ca0",
  2859 => x"00002ca0",
  2860 => x"00002ca8",
  2861 => x"00002ca8",
  2862 => x"00002cb0",
  2863 => x"00002cb0",
  2864 => x"00002cb8",
  2865 => x"00002cb8",
  2866 => x"00002cc0",
  2867 => x"00002cc0",
  2868 => x"00002cc8",
  2869 => x"00002cc8",
  2870 => x"00002cd0",
  2871 => x"00002cd0",
  2872 => x"00002cd8",
  2873 => x"00002cd8",
  2874 => x"00002ce0",
  2875 => x"00002ce0",
  2876 => x"00002ce8",
  2877 => x"00002ce8",
  2878 => x"00002cf0",
  2879 => x"00002cf0",
  2880 => x"00002cf8",
  2881 => x"00002cf8",
  2882 => x"00002d00",
  2883 => x"00002d00",
  2884 => x"00002d08",
  2885 => x"00002d08",
  2886 => x"00002d10",
  2887 => x"00002d10",
  2888 => x"00002d18",
  2889 => x"00002d18",
  2890 => x"00002d20",
  2891 => x"00002d20",
  2892 => x"00002d28",
  2893 => x"00002d28",
  2894 => x"00002d30",
  2895 => x"00002d30",
  2896 => x"00002d38",
  2897 => x"00002d38",
  2898 => x"00002d40",
  2899 => x"00002d40",
  2900 => x"00002d48",
  2901 => x"00002d48",
  2902 => x"00002d50",
  2903 => x"00002d50",
  2904 => x"00002d58",
  2905 => x"00002d58",
  2906 => x"00002d60",
  2907 => x"00002d60",
  2908 => x"00002d68",
  2909 => x"00002d68",
  2910 => x"00002d70",
  2911 => x"00002d70",
  2912 => x"00002d78",
  2913 => x"00002d78",
  2914 => x"00002d80",
  2915 => x"00002d80",
  2916 => x"00002d88",
  2917 => x"00002d88",
  2918 => x"00002d90",
  2919 => x"00002d90",
  2920 => x"00002d98",
  2921 => x"00002d98",
  2922 => x"00002da0",
  2923 => x"00002da0",
  2924 => x"00002da8",
  2925 => x"00002da8",
  2926 => x"00002db0",
  2927 => x"00002db0",
  2928 => x"00002db8",
  2929 => x"00002db8",
  2930 => x"00002dc0",
  2931 => x"00002dc0",
  2932 => x"00002dc8",
  2933 => x"00002dc8",
  2934 => x"00002dd0",
  2935 => x"00002dd0",
  2936 => x"00002dd8",
  2937 => x"00002dd8",
  2938 => x"00002de0",
  2939 => x"00002de0",
  2940 => x"00002de8",
  2941 => x"00002de8",
  2942 => x"00002df0",
  2943 => x"00002df0",
  2944 => x"00002df8",
  2945 => x"00002df8",
  2946 => x"00002e00",
  2947 => x"00002e00",
  2948 => x"00002e08",
  2949 => x"00002e08",
  2950 => x"00002e10",
  2951 => x"00002e10",
  2952 => x"00002e18",
  2953 => x"00002e18",
  2954 => x"00002e20",
  2955 => x"00002e20",
  2956 => x"00002e28",
  2957 => x"00002e28",
  2958 => x"00002e30",
  2959 => x"00002e30",
  2960 => x"00002e38",
  2961 => x"00002e38",
  2962 => x"00002e40",
  2963 => x"00002e40",
  2964 => x"00002e48",
  2965 => x"00002e48",
  2966 => x"00002e50",
  2967 => x"00002e50",
  2968 => x"00002e58",
  2969 => x"00002e58",
  2970 => x"00002e60",
  2971 => x"00002e60",
  2972 => x"00002e68",
  2973 => x"00002e68",
  2974 => x"00002e70",
  2975 => x"00002e70",
  2976 => x"00002e78",
  2977 => x"00002e78",
  2978 => x"00002e80",
  2979 => x"00002e80",
  2980 => x"00002e88",
  2981 => x"00002e88",
  2982 => x"00002e90",
  2983 => x"00002e90",
  2984 => x"00002e98",
  2985 => x"00002e98",
  2986 => x"00002ea0",
  2987 => x"00002ea0",
  2988 => x"00002ea8",
  2989 => x"00002ea8",
  2990 => x"00002eb0",
  2991 => x"00002eb0",
  2992 => x"00002eb8",
  2993 => x"00002eb8",
  2994 => x"00002ec0",
  2995 => x"00002ec0",
  2996 => x"00002ec8",
  2997 => x"00002ec8",
  2998 => x"00002ed0",
  2999 => x"00002ed0",
  3000 => x"00002ed8",
  3001 => x"00002ed8",
  3002 => x"00002ee0",
  3003 => x"00002ee0",
  3004 => x"00002ee8",
  3005 => x"00002ee8",
  3006 => x"00002ef0",
  3007 => x"00002ef0",
  3008 => x"00002ef8",
  3009 => x"00002ef8",
  3010 => x"00002f00",
  3011 => x"00002f00",
  3012 => x"00002f08",
  3013 => x"00002f08",
  3014 => x"00002f10",
  3015 => x"00002f10",
  3016 => x"00002f18",
  3017 => x"00002f18",
  3018 => x"00002f20",
  3019 => x"00002f20",
  3020 => x"00002f28",
  3021 => x"00002f28",
  3022 => x"00002f30",
  3023 => x"00002f30",
  3024 => x"00002f38",
  3025 => x"00002f38",
  3026 => x"00002f40",
  3027 => x"00002f40",
  3028 => x"00002f48",
  3029 => x"00002f48",
  3030 => x"00002f50",
  3031 => x"00002f50",
  3032 => x"00002f58",
  3033 => x"00002f58",
  3034 => x"00002f60",
  3035 => x"00002f60",
  3036 => x"00002f68",
  3037 => x"00002f68",
  3038 => x"00002f70",
  3039 => x"00002f70",
  3040 => x"00002f78",
  3041 => x"00002f78",
  3042 => x"00002f80",
  3043 => x"00002f80",
  3044 => x"00002f88",
  3045 => x"00002f88",
  3046 => x"00002f90",
  3047 => x"00002f90",
  3048 => x"000027b0",
  3049 => x"ffffffff",
  3050 => x"00000000",
  3051 => x"ffffffff",
  3052 => x"00000000",
  3053 => x"00000000",
  others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture rtl; -- Entity: SinglePortRAM

